`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    02:59:20 01/14/2020 
// Design Name: 
// Module Name:    LeftBarrelShifter 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module LeftShifter(A,B,C);

	input [31:0] A;
	input [4:0] B;
	output [31:0] C;
	
	wire [31:0] ST1,ST2,ST3,ST4;
	
	MUX2_1 m1_0 (1'b0, A[0], ST1[0], B[0]);
	MUX2_1 m1_1 (A[0], A[1], ST1[1], B[0]);
	MUX2_1 m1_2 (A[1], A[2], ST1[2], B[0]);
	MUX2_1 m1_3 (A[2], A[3], ST1[3], B[0]);
	MUX2_1 m1_4 (A[3], A[4], ST1[4], B[0]);
	MUX2_1 m1_5 (A[4], A[5], ST1[5], B[0]);
	MUX2_1 m1_6 (A[5], A[6], ST1[6], B[0]);
	MUX2_1 m1_7 (A[6], A[7], ST1[7], B[0]);
	MUX2_1 m1_8 (A[7], A[8], ST1[8], B[0]);
	MUX2_1 m1_9 (A[8], A[9], ST1[9], B[0]);
	MUX2_1 m1_10 (A[9], A[10], ST1[10], B[0]);
	MUX2_1 m1_11 (A[10], A[11], ST1[11], B[0]);
	MUX2_1 m1_12 (A[11], A[12], ST1[12], B[0]);
	MUX2_1 m1_13 (A[12], A[13], ST1[13], B[0]);
	MUX2_1 m1_14 (A[13], A[14], ST1[14], B[0]);
	MUX2_1 m1_15 (A[14], A[15], ST1[15], B[0]);
	MUX2_1 m1_16 (A[15], A[16], ST1[16], B[0]);
	MUX2_1 m1_17 (A[16], A[17], ST1[17], B[0]);
	MUX2_1 m1_18 (A[17], A[18], ST1[18], B[0]);
	MUX2_1 m1_19 (A[18], A[19], ST1[19], B[0]);
	MUX2_1 m1_20 (A[19], A[20], ST1[20], B[0]);
	MUX2_1 m1_21 (A[20], A[21], ST1[21], B[0]);
	MUX2_1 m1_22 (A[21], A[22], ST1[22], B[0]);
	MUX2_1 m1_23 (A[22], A[23], ST1[23], B[0]);
	MUX2_1 m1_24 (A[23], A[24], ST1[24], B[0]);
	MUX2_1 m1_25 (A[24], A[25], ST1[25], B[0]);
	MUX2_1 m1_26 (A[25], A[26], ST1[26], B[0]);
	MUX2_1 m1_27 (A[26], A[27], ST1[27], B[0]);
	MUX2_1 m1_28 (A[27], A[28], ST1[28], B[0]);
	MUX2_1 m1_29 (A[28], A[29], ST1[29], B[0]);
	MUX2_1 m1_30 (A[29], A[30], ST1[30], B[0]);
	MUX2_1 m1_31 (A[30], A[31], ST1[31], B[0]);
	MUX2_1 m2_0 (1'b0, ST1[0], ST2[0], B[1]);
	MUX2_1 m2_1 (1'b0, ST1[1], ST2[1], B[1]);
	MUX2_1 m2_2 (ST1[0], ST1[2], ST2[2], B[1]);
	MUX2_1 m2_3 (ST1[1], ST1[3], ST2[3], B[1]);
	MUX2_1 m2_4 (ST1[2], ST1[4], ST2[4], B[1]);
	MUX2_1 m2_5 (ST1[3], ST1[5], ST2[5], B[1]);
	MUX2_1 m2_6 (ST1[4], ST1[6], ST2[6], B[1]);
	MUX2_1 m2_7 (ST1[5], ST1[7], ST2[7], B[1]);
	MUX2_1 m2_8 (ST1[6], ST1[8], ST2[8], B[1]);
	MUX2_1 m2_9 (ST1[7], ST1[9], ST2[9], B[1]);
	MUX2_1 m2_10 (ST1[8], ST1[10], ST2[10], B[1]);
	MUX2_1 m2_11 (ST1[9], ST1[11], ST2[11], B[1]);
	MUX2_1 m2_12 (ST1[10], ST1[12], ST2[12], B[1]);
	MUX2_1 m2_13 (ST1[11], ST1[13], ST2[13], B[1]);
	MUX2_1 m2_14 (ST1[12], ST1[14], ST2[14], B[1]);
	MUX2_1 m2_15 (ST1[13], ST1[15], ST2[15], B[1]);
	MUX2_1 m2_16 (ST1[14], ST1[16], ST2[16], B[1]);
	MUX2_1 m2_17 (ST1[15], ST1[17], ST2[17], B[1]);
	MUX2_1 m2_18 (ST1[16], ST1[18], ST2[18], B[1]);
	MUX2_1 m2_19 (ST1[17], ST1[19], ST2[19], B[1]);
	MUX2_1 m2_20 (ST1[18], ST1[20], ST2[20], B[1]);
	MUX2_1 m2_21 (ST1[19], ST1[21], ST2[21], B[1]);
	MUX2_1 m2_22 (ST1[20], ST1[22], ST2[22], B[1]);
	MUX2_1 m2_23 (ST1[21], ST1[23], ST2[23], B[1]);
	MUX2_1 m2_24 (ST1[22], ST1[24], ST2[24], B[1]);
	MUX2_1 m2_25 (ST1[23], ST1[25], ST2[25], B[1]);
	MUX2_1 m2_26 (ST1[24], ST1[26], ST2[26], B[1]);
	MUX2_1 m2_27 (ST1[25], ST1[27], ST2[27], B[1]);
	MUX2_1 m2_28 (ST1[26], ST1[28], ST2[28], B[1]);
	MUX2_1 m2_29 (ST1[27], ST1[29], ST2[29], B[1]);
	MUX2_1 m2_30 (ST1[28], ST1[30], ST2[30], B[1]);
	MUX2_1 m2_31 (ST1[29], ST1[31], ST2[31], B[1]);
	MUX2_1 m3_0 (1'b0, ST2[0], ST3[0], B[2]);
	MUX2_1 m3_1 (1'b0, ST2[1], ST3[1], B[2]);
	MUX2_1 m3_2 (1'b0, ST2[2], ST3[2], B[2]);
	MUX2_1 m3_3 (1'b0, ST2[3], ST3[3], B[2]);
	MUX2_1 m3_4 (ST2[0], ST2[4], ST3[4], B[2]);
	MUX2_1 m3_5 (ST2[1], ST2[5], ST3[5], B[2]);
	MUX2_1 m3_6 (ST2[2], ST2[6], ST3[6], B[2]);
	MUX2_1 m3_7 (ST2[3], ST2[7], ST3[7], B[2]);
	MUX2_1 m3_8 (ST2[4], ST2[8], ST3[8], B[2]);
	MUX2_1 m3_9 (ST2[5], ST2[9], ST3[9], B[2]);
	MUX2_1 m3_10 (ST2[6], ST2[10], ST3[10], B[2]);
	MUX2_1 m3_11 (ST2[7], ST2[11], ST3[11], B[2]);
	MUX2_1 m3_12 (ST2[8], ST2[12], ST3[12], B[2]);
	MUX2_1 m3_13 (ST2[9], ST2[13], ST3[13], B[2]);
	MUX2_1 m3_14 (ST2[10], ST2[14], ST3[14], B[2]);
	MUX2_1 m3_15 (ST2[11], ST2[15], ST3[15], B[2]);
	MUX2_1 m3_16 (ST2[12], ST2[16], ST3[16], B[2]);
	MUX2_1 m3_17 (ST2[13], ST2[17], ST3[17], B[2]);
	MUX2_1 m3_18 (ST2[14], ST2[18], ST3[18], B[2]);
	MUX2_1 m3_19 (ST2[15], ST2[19], ST3[19], B[2]);
	MUX2_1 m3_20 (ST2[16], ST2[20], ST3[20], B[2]);
	MUX2_1 m3_21 (ST2[17], ST2[21], ST3[21], B[2]);
	MUX2_1 m3_22 (ST2[18], ST2[22], ST3[22], B[2]);
	MUX2_1 m3_23 (ST2[19], ST2[23], ST3[23], B[2]);
	MUX2_1 m3_24 (ST2[20], ST2[24], ST3[24], B[2]);
	MUX2_1 m3_25 (ST2[21], ST2[25], ST3[25], B[2]);
	MUX2_1 m3_26 (ST2[22], ST2[26], ST3[26], B[2]);
	MUX2_1 m3_27 (ST2[23], ST2[27], ST3[27], B[2]);
	MUX2_1 m3_28 (ST2[24], ST2[28], ST3[28], B[2]);
	MUX2_1 m3_29 (ST2[25], ST2[29], ST3[29], B[2]);
	MUX2_1 m3_30 (ST2[26], ST2[30], ST3[30], B[2]);
	MUX2_1 m3_31 (ST2[27], ST2[31], ST3[31], B[2]);
	MUX2_1 m4_0 (1'b0, ST3[0], ST4[0], B[3]);
	MUX2_1 m4_1 (1'b0, ST3[1], ST4[1], B[3]);
	MUX2_1 m4_2 (1'b0, ST3[2], ST4[2], B[3]);
	MUX2_1 m4_3 (1'b0, ST3[3], ST4[3], B[3]);
	MUX2_1 m4_4 (1'b0, ST3[4], ST4[4], B[3]);
	MUX2_1 m4_5 (1'b0, ST3[5], ST4[5], B[3]);
	MUX2_1 m4_6 (1'b0, ST3[6], ST4[6], B[3]);
	MUX2_1 m4_7 (1'b0, ST3[7], ST4[7], B[3]);
	MUX2_1 m4_8 (ST3[0], ST3[8], ST4[8], B[3]);
	MUX2_1 m4_9 (ST3[1], ST3[9], ST4[9], B[3]);
	MUX2_1 m4_10 (ST3[2], ST3[10], ST4[10], B[3]);
	MUX2_1 m4_11 (ST3[3], ST3[11], ST4[11], B[3]);
	MUX2_1 m4_12 (ST3[4], ST3[12], ST4[12], B[3]);
	MUX2_1 m4_13 (ST3[5], ST3[13], ST4[13], B[3]);
	MUX2_1 m4_14 (ST3[6], ST3[14], ST4[14], B[3]);
	MUX2_1 m4_15 (ST3[7], ST3[15], ST4[15], B[3]);
	MUX2_1 m4_16 (ST3[8], ST3[16], ST4[16], B[3]);
	MUX2_1 m4_17 (ST3[9], ST3[17], ST4[17], B[3]);
	MUX2_1 m4_18 (ST3[10], ST3[18], ST4[18], B[3]);
	MUX2_1 m4_19 (ST3[11], ST3[19], ST4[19], B[3]);
	MUX2_1 m4_20 (ST3[12], ST3[20], ST4[20], B[3]);
	MUX2_1 m4_21 (ST3[13], ST3[21], ST4[21], B[3]);
	MUX2_1 m4_22 (ST3[14], ST3[22], ST4[22], B[3]);
	MUX2_1 m4_23 (ST3[15], ST3[23], ST4[23], B[3]);
	MUX2_1 m4_24 (ST3[16], ST3[24], ST4[24], B[3]);
	MUX2_1 m4_25 (ST3[17], ST3[25], ST4[25], B[3]);
	MUX2_1 m4_26 (ST3[18], ST3[26], ST4[26], B[3]);
	MUX2_1 m4_27 (ST3[19], ST3[27], ST4[27], B[3]);
	MUX2_1 m4_28 (ST3[20], ST3[28], ST4[28], B[3]);
	MUX2_1 m4_29 (ST3[21], ST3[29], ST4[29], B[3]);
	MUX2_1 m4_30 (ST3[22], ST3[30], ST4[30], B[3]);
	MUX2_1 m4_31 (ST3[23], ST3[31], ST4[31], B[3]);
	MUX2_1 m5_0 (1'b0, ST4[0], C[0], B[4]);
	MUX2_1 m5_1 (1'b0, ST4[1], C[1], B[4]);
	MUX2_1 m5_2 (1'b0, ST4[2], C[2], B[4]);
	MUX2_1 m5_3 (1'b0, ST4[3], C[3], B[4]);
	MUX2_1 m5_4 (1'b0, ST4[4], C[4], B[4]);
	MUX2_1 m5_5 (1'b0, ST4[5], C[5], B[4]);
	MUX2_1 m5_6 (1'b0, ST4[6], C[6], B[4]);
	MUX2_1 m5_7 (1'b0, ST4[7], C[7], B[4]);
	MUX2_1 m5_8 (1'b0, ST4[8], C[8], B[4]);
	MUX2_1 m5_9 (1'b0, ST4[9], C[9], B[4]);
	MUX2_1 m5_10 (1'b0, ST4[10], C[10], B[4]);
	MUX2_1 m5_11 (1'b0, ST4[11], C[11], B[4]);
	MUX2_1 m5_12 (1'b0, ST4[12], C[12], B[4]);
	MUX2_1 m5_13 (1'b0, ST4[13], C[13], B[4]);
	MUX2_1 m5_14 (1'b0, ST4[14], C[14], B[4]);
	MUX2_1 m5_15 (1'b0, ST4[15], C[15], B[4]);
	MUX2_1 m5_16 (ST4[0], ST4[16], C[16], B[4]);
	MUX2_1 m5_17 (ST4[1], ST4[17], C[17], B[4]);
	MUX2_1 m5_18 (ST4[2], ST4[18], C[18], B[4]);
	MUX2_1 m5_19 (ST4[3], ST4[19], C[19], B[4]);
	MUX2_1 m5_20 (ST4[4], ST4[20], C[20], B[4]);
	MUX2_1 m5_21 (ST4[5], ST4[21], C[21], B[4]);
	MUX2_1 m5_22 (ST4[6], ST4[22], C[22], B[4]);
	MUX2_1 m5_23 (ST4[7], ST4[23], C[23], B[4]);
	MUX2_1 m5_24 (ST4[8], ST4[24], C[24], B[4]);
	MUX2_1 m5_25 (ST4[9], ST4[25], C[25], B[4]);
	MUX2_1 m5_26 (ST4[10], ST4[26], C[26], B[4]);
	MUX2_1 m5_27 (ST4[11], ST4[27], C[27], B[4]);
	MUX2_1 m5_28 (ST4[12], ST4[28], C[28], B[4]);
	MUX2_1 m5_29 (ST4[13], ST4[29], C[29], B[4]);
	MUX2_1 m5_30 (ST4[14], ST4[30], C[30], B[4]);
	MUX2_1 m5_31 (ST4[15], ST4[31], C[31], B[4]);
endmodule
